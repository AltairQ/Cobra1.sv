// ps2.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module ps2 (
		input  wire       clk_clk,             //                           clk.clk
		input  wire [7:0] ps2_0_command,       // ps2_0_avalon_ps2_command_sink.data
		input  wire       ps2_0_command_valid, //                              .valid
		output wire       ps2_0_command_ready, //                              .ready
		input  wire       ps2_0_data_ready,    //  ps2_0_avalon_ps2_data_source.ready
		output wire [7:0] ps2_0_data,          //                              .data
		output wire       ps2_0_data_valid,    //                              .valid
		inout  wire       ps2_0_PS2_CLK,       //      ps2_0_external_interface.CLK
		inout  wire       ps2_0_PS2_DAT,       //                              .DAT
		input  wire       reset_reset_n        //                         reset.reset_n
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> ps2_0:reset

	ps2_ps2_0 ps2_0 (
		.clk           (clk_clk),                        //                     clk.clk
		.reset         (rst_controller_reset_out_reset), //                   reset.reset
		.command       (ps2_0_command),                  // avalon_ps2_command_sink.data
		.command_valid (ps2_0_command_valid),            //                        .valid
		.command_ready (ps2_0_command_ready),            //                        .ready
		.data_ready    (ps2_0_data_ready),               //  avalon_ps2_data_source.ready
		.data          (ps2_0_data),                     //                        .data
		.data_valid    (ps2_0_data_valid),               //                        .valid
		.PS2_CLK       (ps2_0_PS2_CLK),                  //      external_interface.export
		.PS2_DAT       (ps2_0_PS2_DAT)                   //                        .export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
